module Sprite(
	
	);


endmodule
