module hexaToBinary(
	input [5:0] hexa,
	output [5:0] volteado
	);
	/*
	assign volteado[2]=hexa[0];
	assign volteado[2]=hexa[1];
	
	assign volteado[1]=hexa[1];
	assign volteado[0]=hexa[2];
	*/
	


endmodule 