module WinSpriteCharacter(
	input [9:0] x_pos,y_pos,
	input [9:0] h_count,v_count,
	output logic [23:0] RGB,
	output visible
	);
	logic [9:0] i_pos,j_pos;
	logic [2:0] sprite [0:31][0:31];
	assign sprite= '{
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000, 3'b000}, 
	'{3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000}, 
	'{3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000}, 
	'{3'b000, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b000}, 
	'{3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010}, 
	'{3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010}, 
	'{3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b011, 3'b010, 3'b011, 3'b011, 3'b010, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b100, 3'b010}, 
	'{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b011, 3'b010, 3'b011, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010}, 
	'{3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b001, 3'b011, 3'b010, 3'b011, 3'b011, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010}, 
	'{3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010}, 
	'{3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010}, 
	'{3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010}, 
	'{3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000}, 
	'{3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b010, 3'b010, 3'b010, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000}, 
	'{3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000}, 
	'{3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b001, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b011, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}, 
	'{3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b010, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000, 3'b000}
	};
	
	logic [2:0] codedColor;
	logic inArea;
	spritePositionVerificator spv(x_pos,y_pos,h_count,v_count,inArea,i_pos,j_pos);
	
	assign codedColor=sprite[j_pos][i_pos];
		
		
	//Comparador igual
	logic res [2:0];
	logic S;
	xnor xn1(res[0],codedColor[0],1'b0);
	xnor xn2(res[1],codedColor[1],1'b0);
	xnor xn3(res[2],codedColor[2],1'b0);
	and n1(S,res[0],res[1],res[2]);
	//comparador igual
	
	//dibujar sprite o fondo
	logic notS;
	not comparador(notS,S);
	and and1(visible,notS,inArea);
	//dibujar sprite o fondo
	
	pokeballColorDecoder pokeball(codedColor,RGB);
	

endmodule
